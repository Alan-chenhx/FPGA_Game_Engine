module object3_rom
	(
		input wire clk,
		input wire [6:0] row,
		input wire [3:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [6:0] row_reg;
	reg [3:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @*
	case ({row_reg, col_reg})
		11'b00000000000: color_data = 12'b011011011110;
		11'b00000000001: color_data = 12'b011011011110;
		11'b00000000010: color_data = 12'b011011011110;
		11'b00000000011: color_data = 12'b011011011110;
		11'b00000000100: color_data = 12'b011011011110;
		11'b00000000101: color_data = 12'b011011011110;
		11'b00000000110: color_data = 12'b011011011110;
		11'b00000000111: color_data = 12'b011011011110;
		11'b00000001000: color_data = 12'b011011011110;
		11'b00000001001: color_data = 12'b000000000000;
		11'b00000001010: color_data = 12'b000000000000;
		11'b00000001011: color_data = 12'b011011011110;
		11'b00000001100: color_data = 12'b011011011110;
		11'b00000001101: color_data = 12'b011011011110;
		11'b00000001110: color_data = 12'b011011011110;
		11'b00000001111: color_data = 12'b011011011110;

		11'b00000010000: color_data = 12'b011011011110;
		11'b00000010001: color_data = 12'b011011011110;
		11'b00000010010: color_data = 12'b011011011110;
		11'b00000010011: color_data = 12'b011011011110;
		11'b00000010100: color_data = 12'b011011011110;
		11'b00000010101: color_data = 12'b011011011110;
		11'b00000010110: color_data = 12'b011011011110;
		11'b00000010111: color_data = 12'b011011011110;
		11'b00000011000: color_data = 12'b000000000000;
		11'b00000011001: color_data = 12'b000001110000;
		11'b00000011010: color_data = 12'b000011110000;
		11'b00000011011: color_data = 12'b000000000000;
		11'b00000011100: color_data = 12'b011011011110;
		11'b00000011101: color_data = 12'b011011011110;
		11'b00000011110: color_data = 12'b011011011110;
		11'b00000011111: color_data = 12'b011011011110;

		11'b00000100000: color_data = 12'b011011011110;
		11'b00000100001: color_data = 12'b011011011110;
		11'b00000100010: color_data = 12'b011011011110;
		11'b00000100011: color_data = 12'b011011011110;
		11'b00000100100: color_data = 12'b011011011110;
		11'b00000100101: color_data = 12'b011011011110;
		11'b00000100110: color_data = 12'b011011011110;
		11'b00000100111: color_data = 12'b011011011110;
		11'b00000101000: color_data = 12'b111111111111;
		11'b00000101001: color_data = 12'b111111111111;
		11'b00000101010: color_data = 12'b000001110000;
		11'b00000101011: color_data = 12'b000010110000;
		11'b00000101100: color_data = 12'b000000000000;
		11'b00000101101: color_data = 12'b011011011110;
		11'b00000101110: color_data = 12'b011011011110;
		11'b00000101111: color_data = 12'b011011011110;

		11'b00000110000: color_data = 12'b011011011110;
		11'b00000110001: color_data = 12'b011011011110;
		11'b00000110010: color_data = 12'b011011011110;
		11'b00000110011: color_data = 12'b011011011110;
		11'b00000110100: color_data = 12'b011011011110;
		11'b00000110101: color_data = 12'b011011011110;
		11'b00000110110: color_data = 12'b011011011110;
		11'b00000110111: color_data = 12'b011011011110;
		11'b00000111000: color_data = 12'b000000000000;
		11'b00000111001: color_data = 12'b111111111111;
		11'b00000111010: color_data = 12'b111111111111;
		11'b00000111011: color_data = 12'b000001110000;
		11'b00000111100: color_data = 12'b000000000000;
		11'b00000111101: color_data = 12'b011011011110;
		11'b00000111110: color_data = 12'b011011011110;
		11'b00000111111: color_data = 12'b011011011110;

		11'b00001000000: color_data = 12'b011011011110;
		11'b00001000001: color_data = 12'b011011011110;
		11'b00001000010: color_data = 12'b011011011110;
		11'b00001000011: color_data = 12'b011011011110;
		11'b00001000100: color_data = 12'b000000000000;
		11'b00001000101: color_data = 12'b000000000000;
		11'b00001000110: color_data = 12'b000000000000;
		11'b00001000111: color_data = 12'b011011011110;
		11'b00001001000: color_data = 12'b000000000000;
		11'b00001001001: color_data = 12'b111111111111;
		11'b00001001010: color_data = 12'b111111111111;
		11'b00001001011: color_data = 12'b111111111111;
		11'b00001001100: color_data = 12'b000000000000;
		11'b00001001101: color_data = 12'b000000000000;
		11'b00001001110: color_data = 12'b000000000000;
		11'b00001001111: color_data = 12'b011011011110;

		11'b00001010000: color_data = 12'b011011011110;
		11'b00001010001: color_data = 12'b011011011110;
		11'b00001010010: color_data = 12'b000000000000;
		11'b00001010011: color_data = 12'b000000000000;
		11'b00001010100: color_data = 12'b000011110000;
		11'b00001010101: color_data = 12'b000011110000;
		11'b00001010110: color_data = 12'b000011110000;
		11'b00001010111: color_data = 12'b000000000000;
		11'b00001011000: color_data = 12'b111111111111;
		11'b00001011001: color_data = 12'b111111111111;
		11'b00001011010: color_data = 12'b111111111111;
		11'b00001011011: color_data = 12'b111111111111;
		11'b00001011100: color_data = 12'b000000000000;
		11'b00001011101: color_data = 12'b111110000000;
		11'b00001011110: color_data = 12'b111110000000;
		11'b00001011111: color_data = 12'b000000000000;

		11'b00001100000: color_data = 12'b011011011110;
		11'b00001100001: color_data = 12'b000000000000;
		11'b00001100010: color_data = 12'b000011110000;
		11'b00001100011: color_data = 12'b111111111111;
		11'b00001100100: color_data = 12'b111111111111;
		11'b00001100101: color_data = 12'b000011110000;
		11'b00001100110: color_data = 12'b000011110000;
		11'b00001100111: color_data = 12'b000011110000;
		11'b00001101000: color_data = 12'b000001110000;
		11'b00001101001: color_data = 12'b111111111111;
		11'b00001101010: color_data = 12'b111111111111;
		11'b00001101011: color_data = 12'b000001110000;
		11'b00001101100: color_data = 12'b000000000000;
		11'b00001101101: color_data = 12'b111110000000;
		11'b00001101110: color_data = 12'b111110000000;
		11'b00001101111: color_data = 12'b000000000000;

		11'b00001110000: color_data = 12'b011011011110;
		11'b00001110001: color_data = 12'b000000000000;
		11'b00001110010: color_data = 12'b111111111111;
		11'b00001110011: color_data = 12'b000000000000;
		11'b00001110100: color_data = 12'b000011110000;
		11'b00001110101: color_data = 12'b000011110000;
		11'b00001110110: color_data = 12'b000011110000;
		11'b00001110111: color_data = 12'b000011110000;
		11'b00001111000: color_data = 12'b000011110000;
		11'b00001111001: color_data = 12'b000001110000;
		11'b00001111010: color_data = 12'b000001110000;
		11'b00001111011: color_data = 12'b000010110000;
		11'b00001111100: color_data = 12'b000000000000;
		11'b00001111101: color_data = 12'b000000000000;
		11'b00001111110: color_data = 12'b000000000000;
		11'b00001111111: color_data = 12'b011011011110;

		11'b00010000000: color_data = 12'b000000000000;
		11'b00010000001: color_data = 12'b000011110000;
		11'b00010000010: color_data = 12'b000011110000;
		11'b00010000011: color_data = 12'b000011110000;
		11'b00010000100: color_data = 12'b000011110000;
		11'b00010000101: color_data = 12'b000011110000;
		11'b00010000110: color_data = 12'b000011110000;
		11'b00010000111: color_data = 12'b000011110000;
		11'b00010001000: color_data = 12'b000011110000;
		11'b00010001001: color_data = 12'b000011110000;
		11'b00010001010: color_data = 12'b000010110000;
		11'b00010001011: color_data = 12'b000010110000;
		11'b00010001100: color_data = 12'b000001110000;
		11'b00010001101: color_data = 12'b000000000000;
		11'b00010001110: color_data = 12'b111110000000;
		11'b00010001111: color_data = 12'b000000000000;

		11'b00010010000: color_data = 12'b000000000000;
		11'b00010010001: color_data = 12'b000011110000;
		11'b00010010010: color_data = 12'b000011110000;
		11'b00010010011: color_data = 12'b000011110000;
		11'b00010010100: color_data = 12'b000011110000;
		11'b00010010101: color_data = 12'b000011110000;
		11'b00010010110: color_data = 12'b000010110000;
		11'b00010010111: color_data = 12'b000011110000;
		11'b00010011000: color_data = 12'b000011110000;
		11'b00010011001: color_data = 12'b000011110000;
		11'b00010011010: color_data = 12'b000011110000;
		11'b00010011011: color_data = 12'b000010110000;
		11'b00010011100: color_data = 12'b000001110000;
		11'b00010011101: color_data = 12'b000000000000;
		11'b00010011110: color_data = 12'b111110000000;
		11'b00010011111: color_data = 12'b000000000000;

		11'b00010100000: color_data = 12'b000000000000;
		11'b00010100001: color_data = 12'b000011110000;
		11'b00010100010: color_data = 12'b000011110000;
		11'b00010100011: color_data = 12'b000011110000;
		11'b00010100100: color_data = 12'b000011110000;
		11'b00010100101: color_data = 12'b000010110000;
		11'b00010100110: color_data = 12'b000000000000;
		11'b00010100111: color_data = 12'b111111111111;
		11'b00010101000: color_data = 12'b000011110000;
		11'b00010101001: color_data = 12'b000011110000;
		11'b00010101010: color_data = 12'b000011110000;
		11'b00010101011: color_data = 12'b000010110000;
		11'b00010101100: color_data = 12'b000001110000;
		11'b00010101101: color_data = 12'b000000000000;
		11'b00010101110: color_data = 12'b000000000000;
		11'b00010101111: color_data = 12'b011011011110;

		11'b00010110000: color_data = 12'b000000000000;
		11'b00010110001: color_data = 12'b000011110000;
		11'b00010110010: color_data = 12'b000011110000;
		11'b00010110011: color_data = 12'b000011110000;
		11'b00010110100: color_data = 12'b000011110000;
		11'b00010110101: color_data = 12'b000010110000;
		11'b00010110110: color_data = 12'b000000000000;
		11'b00010110111: color_data = 12'b111111111111;
		11'b00010111000: color_data = 12'b000011110000;
		11'b00010111001: color_data = 12'b000011110000;
		11'b00010111010: color_data = 12'b000011110000;
		11'b00010111011: color_data = 12'b000010110000;
		11'b00010111100: color_data = 12'b000000000000;
		11'b00010111101: color_data = 12'b111110000000;
		11'b00010111110: color_data = 12'b000000000000;
		11'b00010111111: color_data = 12'b011011011110;

		11'b00011000000: color_data = 12'b000000000000;
		11'b00011000001: color_data = 12'b000010110000;
		11'b00011000010: color_data = 12'b000011110000;
		11'b00011000011: color_data = 12'b000011110000;
		11'b00011000100: color_data = 12'b000010110000;
		11'b00011000101: color_data = 12'b000001110000;
		11'b00011000110: color_data = 12'b000000000000;
		11'b00011000111: color_data = 12'b000000000000;
		11'b00011001000: color_data = 12'b111111111111;
		11'b00011001001: color_data = 12'b000011110000;
		11'b00011001010: color_data = 12'b000011110000;
		11'b00011001011: color_data = 12'b000010110000;
		11'b00011001100: color_data = 12'b000000000000;
		11'b00011001101: color_data = 12'b111110000000;
		11'b00011001110: color_data = 12'b000000000000;
		11'b00011001111: color_data = 12'b011011011110;

		11'b00011010000: color_data = 12'b011011011110;
		11'b00011010001: color_data = 12'b000000000000;
		11'b00011010010: color_data = 12'b000010110000;
		11'b00011010011: color_data = 12'b000010110000;
		11'b00011010100: color_data = 12'b000001110000;
		11'b00011010101: color_data = 12'b000000000000;
		11'b00011010110: color_data = 12'b111111111111;
		11'b00011010111: color_data = 12'b111111111111;
		11'b00011011000: color_data = 12'b111111111111;
		11'b00011011001: color_data = 12'b111111111111;
		11'b00011011010: color_data = 12'b111111111111;
		11'b00011011011: color_data = 12'b000010110000;
		11'b00011011100: color_data = 12'b000000000000;
		11'b00011011101: color_data = 12'b000000000000;
		11'b00011011110: color_data = 12'b000000000000;
		11'b00011011111: color_data = 12'b011011011110;

		11'b00011100000: color_data = 12'b011011011110;
		11'b00011100001: color_data = 12'b011011011110;
		11'b00011100010: color_data = 12'b000000000000;
		11'b00011100011: color_data = 12'b000000000000;
		11'b00011100100: color_data = 12'b000000000000;
		11'b00011100101: color_data = 12'b111111111111;
		11'b00011100110: color_data = 12'b111111111111;
		11'b00011100111: color_data = 12'b111111111111;
		11'b00011101000: color_data = 12'b000000000000;
		11'b00011101001: color_data = 12'b111111111111;
		11'b00011101010: color_data = 12'b111111111111;
		11'b00011101011: color_data = 12'b000010110000;
		11'b00011101100: color_data = 12'b000001110000;
		11'b00011101101: color_data = 12'b000000000000;
		11'b00011101110: color_data = 12'b111110000000;
		11'b00011101111: color_data = 12'b000000000000;

		11'b00011110000: color_data = 12'b011011011110;
		11'b00011110001: color_data = 12'b011011011110;
		11'b00011110010: color_data = 12'b011011011110;
		11'b00011110011: color_data = 12'b011011011110;
		11'b00011110100: color_data = 12'b011011011110;
		11'b00011110101: color_data = 12'b000000000000;
		11'b00011110110: color_data = 12'b000000000000;
		11'b00011110111: color_data = 12'b000000000000;
		11'b00011111000: color_data = 12'b011011011110;
		11'b00011111001: color_data = 12'b000000000000;
		11'b00011111010: color_data = 12'b111111111111;
		11'b00011111011: color_data = 12'b000010110000;
		11'b00011111100: color_data = 12'b000010110000;
		11'b00011111101: color_data = 12'b000000000000;
		11'b00011111110: color_data = 12'b000000000000;
		11'b00011111111: color_data = 12'b011011011110;

		11'b00100000000: color_data = 12'b000000000000;
		11'b00100000001: color_data = 12'b111111111111;
		11'b00100000010: color_data = 12'b000010110000;
		11'b00100000011: color_data = 12'b000001110000;
		11'b00100000100: color_data = 12'b000000000000;
		11'b00100000101: color_data = 12'b000000000000;
		11'b00100000110: color_data = 12'b011011011110;
		11'b00100000111: color_data = 12'b000000000000;
		11'b00100001000: color_data = 12'b000000000000;
		11'b00100001001: color_data = 12'b000000000000;
		11'b00100001010: color_data = 12'b000000000000;
		11'b00100001011: color_data = 12'b011011011110;
		11'b00100001100: color_data = 12'b000000000000;
		11'b00100001101: color_data = 12'b000000000000;
		11'b00100001110: color_data = 12'b011011011110;
		11'b00100001111: color_data = 12'b011011011110;

		11'b00100010000: color_data = 12'b000000000000;
		11'b00100010001: color_data = 12'b111111111111;
		11'b00100010010: color_data = 12'b000011110000;
		11'b00100010011: color_data = 12'b000010110000;
		11'b00100010100: color_data = 12'b000000000000;
		11'b00100010101: color_data = 12'b111111111111;
		11'b00100010110: color_data = 12'b000000000000;
		11'b00100010111: color_data = 12'b111111111111;
		11'b00100011000: color_data = 12'b111110000000;
		11'b00100011001: color_data = 12'b111110000000;
		11'b00100011010: color_data = 12'b101100100000;
		11'b00100011011: color_data = 12'b000000000000;
		11'b00100011100: color_data = 12'b111111111111;
		11'b00100011101: color_data = 12'b000000000000;
		11'b00100011110: color_data = 12'b000000000000;
		11'b00100011111: color_data = 12'b000000000000;

		11'b00100100000: color_data = 12'b000000000000;
		11'b00100100001: color_data = 12'b111111111111;
		11'b00100100010: color_data = 12'b000011110000;
		11'b00100100011: color_data = 12'b000010110000;
		11'b00100100100: color_data = 12'b000000000000;
		11'b00100100101: color_data = 12'b111111111111;
		11'b00100100110: color_data = 12'b000000000000;
		11'b00100100111: color_data = 12'b111110000000;
		11'b00100101000: color_data = 12'b101100100000;
		11'b00100101001: color_data = 12'b101100100000;
		11'b00100101010: color_data = 12'b101100100000;
		11'b00100101011: color_data = 12'b000000000000;
		11'b00100101100: color_data = 12'b111111111111;
		11'b00100101101: color_data = 12'b000000000000;
		11'b00100101110: color_data = 12'b000010110000;
		11'b00100101111: color_data = 12'b000000000000;

		11'b00100110000: color_data = 12'b000000000000;
		11'b00100110001: color_data = 12'b111111111111;
		11'b00100110010: color_data = 12'b111111111111;
		11'b00100110011: color_data = 12'b000011110000;
		11'b00100110100: color_data = 12'b000010110000;
		11'b00100110101: color_data = 12'b000000000000;
		11'b00100110110: color_data = 12'b111111111111;
		11'b00100110111: color_data = 12'b000000000000;
		11'b00100111000: color_data = 12'b000000000000;
		11'b00100111001: color_data = 12'b000000000000;
		11'b00100111010: color_data = 12'b000000000000;
		11'b00100111011: color_data = 12'b111111111111;
		11'b00100111100: color_data = 12'b000000000000;
		11'b00100111101: color_data = 12'b000010110000;
		11'b00100111110: color_data = 12'b000000000000;
		11'b00100111111: color_data = 12'b011011011110;

		11'b00101000000: color_data = 12'b011011011110;
		11'b00101000001: color_data = 12'b000000000000;
		11'b00101000010: color_data = 12'b111111111111;
		11'b00101000011: color_data = 12'b000011110000;
		11'b00101000100: color_data = 12'b000000000000;
		11'b00101000101: color_data = 12'b000000000000;
		11'b00101000110: color_data = 12'b000000000000;
		11'b00101000111: color_data = 12'b111111111111;
		11'b00101001000: color_data = 12'b111111111111;
		11'b00101001001: color_data = 12'b111111111111;
		11'b00101001010: color_data = 12'b111111111111;
		11'b00101001011: color_data = 12'b111111111111;
		11'b00101001100: color_data = 12'b000000000000;
		11'b00101001101: color_data = 12'b000010110000;
		11'b00101001110: color_data = 12'b000000000000;
		11'b00101001111: color_data = 12'b011011011110;

		11'b00101010000: color_data = 12'b011011011110;
		11'b00101010001: color_data = 12'b000000000000;
		11'b00101010010: color_data = 12'b111111111111;
		11'b00101010011: color_data = 12'b000011110000;
		11'b00101010100: color_data = 12'b000000000000;
		11'b00101010101: color_data = 12'b111110000000;
		11'b00101010110: color_data = 12'b111110000000;
		11'b00101010111: color_data = 12'b000000000000;
		11'b00101011000: color_data = 12'b000000000000;
		11'b00101011001: color_data = 12'b000000000000;
		11'b00101011010: color_data = 12'b000000000000;
		11'b00101011011: color_data = 12'b000000000000;
		11'b00101011100: color_data = 12'b000010110000;
		11'b00101011101: color_data = 12'b111111111111;
		11'b00101011110: color_data = 12'b000000000000;
		11'b00101011111: color_data = 12'b011011011110;

		11'b00101100000: color_data = 12'b011011011110;
		11'b00101100001: color_data = 12'b000000000000;
		11'b00101100010: color_data = 12'b111111111111;
		11'b00101100011: color_data = 12'b111111111111;
		11'b00101100100: color_data = 12'b111111111111;
		11'b00101100101: color_data = 12'b000000000000;
		11'b00101100110: color_data = 12'b111110000000;
		11'b00101100111: color_data = 12'b111110000000;
		11'b00101101000: color_data = 12'b000000000000;
		11'b00101101001: color_data = 12'b000010110000;
		11'b00101101010: color_data = 12'b000010110000;
		11'b00101101011: color_data = 12'b000010110000;
		11'b00101101100: color_data = 12'b111111111111;
		11'b00101101101: color_data = 12'b000000000000;
		11'b00101101110: color_data = 12'b011011011110;
		11'b00101101111: color_data = 12'b011011011110;

		11'b00101110000: color_data = 12'b011011011110;
		11'b00101110001: color_data = 12'b011011011110;
		11'b00101110010: color_data = 12'b000000000000;
		11'b00101110011: color_data = 12'b111111111111;
		11'b00101110100: color_data = 12'b111111111111;
		11'b00101110101: color_data = 12'b111111111111;
		11'b00101110110: color_data = 12'b000000000000;
		11'b00101110111: color_data = 12'b111110000000;
		11'b00101111000: color_data = 12'b000000000000;
		11'b00101111001: color_data = 12'b111111111111;
		11'b00101111010: color_data = 12'b111111111111;
		11'b00101111011: color_data = 12'b111111111111;
		11'b00101111100: color_data = 12'b111111111111;
		11'b00101111101: color_data = 12'b000000000000;
		11'b00101111110: color_data = 12'b011011011110;
		11'b00101111111: color_data = 12'b011011011110;

		11'b00110000000: color_data = 12'b011011011110;
		11'b00110000001: color_data = 12'b011011011110;
		11'b00110000010: color_data = 12'b000000000000;
		11'b00110000011: color_data = 12'b111111111111;
		11'b00110000100: color_data = 12'b111111111111;
		11'b00110000101: color_data = 12'b000000000000;
		11'b00110000110: color_data = 12'b111110000000;
		11'b00110000111: color_data = 12'b111110000000;
		11'b00110001000: color_data = 12'b111110000000;
		11'b00110001001: color_data = 12'b000000000000;
		11'b00110001010: color_data = 12'b111111111111;
		11'b00110001011: color_data = 12'b111111111111;
		11'b00110001100: color_data = 12'b000000000000;
		11'b00110001101: color_data = 12'b011011011110;
		11'b00110001110: color_data = 12'b011011011110;
		11'b00110001111: color_data = 12'b011011011110;

		11'b00110010000: color_data = 12'b011011011110;
		11'b00110010001: color_data = 12'b011011011110;
		11'b00110010010: color_data = 12'b011011011110;
		11'b00110010011: color_data = 12'b000000000000;
		11'b00110010100: color_data = 12'b111111111111;
		11'b00110010101: color_data = 12'b000000000000;
		11'b00110010110: color_data = 12'b111110000000;
		11'b00110010111: color_data = 12'b111110000000;
		11'b00110011000: color_data = 12'b111110000000;
		11'b00110011001: color_data = 12'b000000000000;
		11'b00110011010: color_data = 12'b000000000000;
		11'b00110011011: color_data = 12'b111111111111;
		11'b00110011100: color_data = 12'b000000000000;
		11'b00110011101: color_data = 12'b011011011110;
		11'b00110011110: color_data = 12'b011011011110;
		11'b00110011111: color_data = 12'b011011011110;

		11'b00110100000: color_data = 12'b011011011110;
		11'b00110100001: color_data = 12'b011011011110;
		11'b00110100010: color_data = 12'b011011011110;
		11'b00110100011: color_data = 12'b011011011110;
		11'b00110100100: color_data = 12'b000000000000;
		11'b00110100101: color_data = 12'b111111111111;
		11'b00110100110: color_data = 12'b000000000000;
		11'b00110100111: color_data = 12'b000000000000;
		11'b00110101000: color_data = 12'b000000000000;
		11'b00110101001: color_data = 12'b111111111111;
		11'b00110101010: color_data = 12'b000000000000;
		11'b00110101011: color_data = 12'b000000000000;
		11'b00110101100: color_data = 12'b011011011110;
		11'b00110101101: color_data = 12'b011011011110;
		11'b00110101110: color_data = 12'b011011011110;
		11'b00110101111: color_data = 12'b011011011110;

		11'b00110110000: color_data = 12'b011011011110;
		11'b00110110001: color_data = 12'b011011011110;
		11'b00110110010: color_data = 12'b011011011110;
		11'b00110110011: color_data = 12'b011011011110;
		11'b00110110100: color_data = 12'b011011011110;
		11'b00110110101: color_data = 12'b000000000000;
		11'b00110110110: color_data = 12'b000000000000;
		11'b00110110111: color_data = 12'b000000000000;
		11'b00110111000: color_data = 12'b000000000000;
		11'b00110111001: color_data = 12'b000000000000;
		11'b00110111010: color_data = 12'b000000000000;
		11'b00110111011: color_data = 12'b011011011110;
		11'b00110111100: color_data = 12'b011011011110;
		11'b00110111101: color_data = 12'b011011011110;
		11'b00110111110: color_data = 12'b011011011110;
		11'b00110111111: color_data = 12'b011011011110;

		11'b00111000000: color_data = 12'b011011011110;
		11'b00111000001: color_data = 12'b011011011110;
		11'b00111000010: color_data = 12'b011011011110;
		11'b00111000011: color_data = 12'b011011011110;
		11'b00111000100: color_data = 12'b011011011110;
		11'b00111000101: color_data = 12'b000000000000;
		11'b00111000110: color_data = 12'b101100100000;
		11'b00111000111: color_data = 12'b101100100000;
		11'b00111001000: color_data = 12'b101100100000;
		11'b00111001001: color_data = 12'b101100100000;
		11'b00111001010: color_data = 12'b101100100000;
		11'b00111001011: color_data = 12'b000000000000;
		11'b00111001100: color_data = 12'b011011011110;
		11'b00111001101: color_data = 12'b011011011110;
		11'b00111001110: color_data = 12'b011011011110;
		11'b00111001111: color_data = 12'b011011011110;

		11'b00111010000: color_data = 12'b011011011110;
		11'b00111010001: color_data = 12'b011011011110;
		11'b00111010010: color_data = 12'b011011011110;
		11'b00111010011: color_data = 12'b011011011110;
		11'b00111010100: color_data = 12'b000000000000;
		11'b00111010101: color_data = 12'b111111111111;
		11'b00111010110: color_data = 12'b101100100000;
		11'b00111010111: color_data = 12'b101100100000;
		11'b00111011000: color_data = 12'b101100100000;
		11'b00111011001: color_data = 12'b101100100000;
		11'b00111011010: color_data = 12'b101100100000;
		11'b00111011011: color_data = 12'b000000000000;
		11'b00111011100: color_data = 12'b011011011110;
		11'b00111011101: color_data = 12'b011011011110;
		11'b00111011110: color_data = 12'b011011011110;
		11'b00111011111: color_data = 12'b011011011110;

		11'b00111100000: color_data = 12'b011011011110;
		11'b00111100001: color_data = 12'b011011011110;
		11'b00111100010: color_data = 12'b011011011110;
		11'b00111100011: color_data = 12'b011011011110;
		11'b00111100100: color_data = 12'b000000000000;
		11'b00111100101: color_data = 12'b101100100000;
		11'b00111100110: color_data = 12'b101100100000;
		11'b00111100111: color_data = 12'b101100100000;
		11'b00111101000: color_data = 12'b101100100000;
		11'b00111101001: color_data = 12'b101100100000;
		11'b00111101010: color_data = 12'b101100100000;
		11'b00111101011: color_data = 12'b000000000000;
		11'b00111101100: color_data = 12'b011011011110;
		11'b00111101101: color_data = 12'b011011011110;
		11'b00111101110: color_data = 12'b011011011110;
		11'b00111101111: color_data = 12'b011011011110;

		11'b00111110000: color_data = 12'b011011011110;
		11'b00111110001: color_data = 12'b011011011110;
		11'b00111110010: color_data = 12'b011011011110;
		11'b00111110011: color_data = 12'b011011011110;
		11'b00111110100: color_data = 12'b000000000000;
		11'b00111110101: color_data = 12'b000000000000;
		11'b00111110110: color_data = 12'b000000000000;
		11'b00111110111: color_data = 12'b000000000000;
		11'b00111111000: color_data = 12'b000000000000;
		11'b00111111001: color_data = 12'b000000000000;
		11'b00111111010: color_data = 12'b000000000000;
		11'b00111111011: color_data = 12'b000000000000;
		11'b00111111100: color_data = 12'b011011011110;
		11'b00111111101: color_data = 12'b011011011110;
		11'b00111111110: color_data = 12'b011011011110;
		11'b00111111111: color_data = 12'b011011011110;

		11'b01000000000: color_data = 12'b000000000000;
		11'b01000000001: color_data = 12'b111111111111;
		11'b01000000010: color_data = 12'b000010110000;
		11'b01000000011: color_data = 12'b000001110000;
		11'b01000000100: color_data = 12'b000000000000;
		11'b01000000101: color_data = 12'b000000000000;
		11'b01000000110: color_data = 12'b011011011110;
		11'b01000000111: color_data = 12'b000000000000;
		11'b01000001000: color_data = 12'b000000000000;
		11'b01000001001: color_data = 12'b000000000000;
		11'b01000001010: color_data = 12'b000000000000;
		11'b01000001011: color_data = 12'b011011011110;
		11'b01000001100: color_data = 12'b000000000000;
		11'b01000001101: color_data = 12'b000000000000;
		11'b01000001110: color_data = 12'b011011011110;
		11'b01000001111: color_data = 12'b011011011110;

		11'b01000010000: color_data = 12'b000000000000;
		11'b01000010001: color_data = 12'b111111111111;
		11'b01000010010: color_data = 12'b000011110000;
		11'b01000010011: color_data = 12'b000010110000;
		11'b01000010100: color_data = 12'b000000000000;
		11'b01000010101: color_data = 12'b111111111111;
		11'b01000010110: color_data = 12'b000000000000;
		11'b01000010111: color_data = 12'b111111111111;
		11'b01000011000: color_data = 12'b111110000000;
		11'b01000011001: color_data = 12'b111110000000;
		11'b01000011010: color_data = 12'b101100100000;
		11'b01000011011: color_data = 12'b000000000000;
		11'b01000011100: color_data = 12'b111111111111;
		11'b01000011101: color_data = 12'b000000000000;
		11'b01000011110: color_data = 12'b000000000000;
		11'b01000011111: color_data = 12'b000000000000;

		11'b01000100000: color_data = 12'b000000000000;
		11'b01000100001: color_data = 12'b111111111111;
		11'b01000100010: color_data = 12'b000011110000;
		11'b01000100011: color_data = 12'b000010110000;
		11'b01000100100: color_data = 12'b000000000000;
		11'b01000100101: color_data = 12'b111111111111;
		11'b01000100110: color_data = 12'b000000000000;
		11'b01000100111: color_data = 12'b111110000000;
		11'b01000101000: color_data = 12'b101100100000;
		11'b01000101001: color_data = 12'b101100100000;
		11'b01000101010: color_data = 12'b101100100000;
		11'b01000101011: color_data = 12'b000000000000;
		11'b01000101100: color_data = 12'b111111111111;
		11'b01000101101: color_data = 12'b000000000000;
		11'b01000101110: color_data = 12'b000010110000;
		11'b01000101111: color_data = 12'b000000000000;

		11'b01000110000: color_data = 12'b000000000000;
		11'b01000110001: color_data = 12'b111111111111;
		11'b01000110010: color_data = 12'b000011110000;
		11'b01000110011: color_data = 12'b000010110000;
		11'b01000110100: color_data = 12'b000010110000;
		11'b01000110101: color_data = 12'b000000000000;
		11'b01000110110: color_data = 12'b111111111111;
		11'b01000110111: color_data = 12'b000000000000;
		11'b01000111000: color_data = 12'b000000000000;
		11'b01000111001: color_data = 12'b000000000000;
		11'b01000111010: color_data = 12'b000000000000;
		11'b01000111011: color_data = 12'b111111111111;
		11'b01000111100: color_data = 12'b000000000000;
		11'b01000111101: color_data = 12'b000010110000;
		11'b01000111110: color_data = 12'b000000000000;
		11'b01000111111: color_data = 12'b011011011110;

		11'b01001000000: color_data = 12'b000000000000;
		11'b01001000001: color_data = 12'b111111111111;
		11'b01001000010: color_data = 12'b111111111111;
		11'b01001000011: color_data = 12'b000011110000;
		11'b01001000100: color_data = 12'b000000000000;
		11'b01001000101: color_data = 12'b111110000000;
		11'b01001000110: color_data = 12'b000000000000;
		11'b01001000111: color_data = 12'b111111111111;
		11'b01001001000: color_data = 12'b111111111111;
		11'b01001001001: color_data = 12'b111111111111;
		11'b01001001010: color_data = 12'b111111111111;
		11'b01001001011: color_data = 12'b111111111111;
		11'b01001001100: color_data = 12'b000000000000;
		11'b01001001101: color_data = 12'b000010110000;
		11'b01001001110: color_data = 12'b000000000000;
		11'b01001001111: color_data = 12'b011011011110;

		11'b01001010000: color_data = 12'b000000000000;
		11'b01001010001: color_data = 12'b111111111111;
		11'b01001010010: color_data = 12'b000000000000;
		11'b01001010011: color_data = 12'b000000000000;
		11'b01001010100: color_data = 12'b000000000000;
		11'b01001010101: color_data = 12'b111110000000;
		11'b01001010110: color_data = 12'b000000000000;
		11'b01001010111: color_data = 12'b000000000000;
		11'b01001011000: color_data = 12'b000000000000;
		11'b01001011001: color_data = 12'b000000000000;
		11'b01001011010: color_data = 12'b000000000000;
		11'b01001011011: color_data = 12'b000000000000;
		11'b01001011100: color_data = 12'b000010110000;
		11'b01001011101: color_data = 12'b111111111111;
		11'b01001011110: color_data = 12'b000000000000;
		11'b01001011111: color_data = 12'b011011011110;

		11'b01001100000: color_data = 12'b011011011110;
		11'b01001100001: color_data = 12'b000000000000;
		11'b01001100010: color_data = 12'b111110000000;
		11'b01001100011: color_data = 12'b111110000000;
		11'b01001100100: color_data = 12'b000000000000;
		11'b01001100101: color_data = 12'b111110000000;
		11'b01001100110: color_data = 12'b000000000000;
		11'b01001100111: color_data = 12'b000010110000;
		11'b01001101000: color_data = 12'b000010110000;
		11'b01001101001: color_data = 12'b000010110000;
		11'b01001101010: color_data = 12'b000010110000;
		11'b01001101011: color_data = 12'b000010110000;
		11'b01001101100: color_data = 12'b111111111111;
		11'b01001101101: color_data = 12'b000000000000;
		11'b01001101110: color_data = 12'b011011011110;
		11'b01001101111: color_data = 12'b011011011110;

		11'b01001110000: color_data = 12'b011011011110;
		11'b01001110001: color_data = 12'b000000000000;
		11'b01001110010: color_data = 12'b111110000000;
		11'b01001110011: color_data = 12'b111110000000;
		11'b01001110100: color_data = 12'b111110000000;
		11'b01001110101: color_data = 12'b111110000000;
		11'b01001110110: color_data = 12'b000000000000;
		11'b01001110111: color_data = 12'b111111111111;
		11'b01001111000: color_data = 12'b000000000000;
		11'b01001111001: color_data = 12'b000000000000;
		11'b01001111010: color_data = 12'b111111111111;
		11'b01001111011: color_data = 12'b111111111111;
		11'b01001111100: color_data = 12'b111111111111;
		11'b01001111101: color_data = 12'b000000000000;
		11'b01001111110: color_data = 12'b011011011110;
		11'b01001111111: color_data = 12'b011011011110;

		11'b01010000000: color_data = 12'b011011011110;
		11'b01010000001: color_data = 12'b011011011110;
		11'b01010000010: color_data = 12'b000000000000;
		11'b01010000011: color_data = 12'b111110000000;
		11'b01010000100: color_data = 12'b111110000000;
		11'b01010000101: color_data = 12'b000000000000;
		11'b01010000110: color_data = 12'b111111111111;
		11'b01010000111: color_data = 12'b000000000000;
		11'b01010001000: color_data = 12'b000010110000;
		11'b01010001001: color_data = 12'b000011110000;
		11'b01010001010: color_data = 12'b000000000000;
		11'b01010001011: color_data = 12'b000000000000;
		11'b01010001100: color_data = 12'b000000000000;
		11'b01010001101: color_data = 12'b011011011110;
		11'b01010001110: color_data = 12'b011011011110;
		11'b01010001111: color_data = 12'b011011011110;

		11'b01010010000: color_data = 12'b011011011110;
		11'b01010010001: color_data = 12'b011011011110;
		11'b01010010010: color_data = 12'b011011011110;
		11'b01010010011: color_data = 12'b000000000000;
		11'b01010010100: color_data = 12'b000000000000;
		11'b01010010101: color_data = 12'b111111111111;
		11'b01010010110: color_data = 12'b111111111111;
		11'b01010010111: color_data = 12'b000000000000;
		11'b01010011000: color_data = 12'b000010110000;
		11'b01010011001: color_data = 12'b000000000000;
		11'b01010011010: color_data = 12'b101100100000;
		11'b01010011011: color_data = 12'b101100100000;
		11'b01010011100: color_data = 12'b000000000000;
		11'b01010011101: color_data = 12'b011011011110;
		11'b01010011110: color_data = 12'b011011011110;
		11'b01010011111: color_data = 12'b011011011110;

		11'b01010100000: color_data = 12'b011011011110;
		11'b01010100001: color_data = 12'b011011011110;
		11'b01010100010: color_data = 12'b000000000000;
		11'b01010100011: color_data = 12'b000000000000;
		11'b01010100100: color_data = 12'b000000000000;
		11'b01010100101: color_data = 12'b111111111111;
		11'b01010100110: color_data = 12'b111111111111;
		11'b01010100111: color_data = 12'b000000000000;
		11'b01010101000: color_data = 12'b000000000000;
		11'b01010101001: color_data = 12'b101100100000;
		11'b01010101010: color_data = 12'b101100100000;
		11'b01010101011: color_data = 12'b101100100000;
		11'b01010101100: color_data = 12'b101100100000;
		11'b01010101101: color_data = 12'b000000000000;
		11'b01010101110: color_data = 12'b011011011110;
		11'b01010101111: color_data = 12'b011011011110;

		11'b01010110000: color_data = 12'b011011011110;
		11'b01010110001: color_data = 12'b000000000000;
		11'b01010110010: color_data = 12'b111111111111;
		11'b01010110011: color_data = 12'b101100100000;
		11'b01010110100: color_data = 12'b101100100000;
		11'b01010110101: color_data = 12'b000000000000;
		11'b01010110110: color_data = 12'b000000000000;
		11'b01010110111: color_data = 12'b000000000000;
		11'b01010111000: color_data = 12'b101100100000;
		11'b01010111001: color_data = 12'b101100100000;
		11'b01010111010: color_data = 12'b101100100000;
		11'b01010111011: color_data = 12'b101100100000;
		11'b01010111100: color_data = 12'b101100100000;
		11'b01010111101: color_data = 12'b000000000000;
		11'b01010111110: color_data = 12'b011011011110;
		11'b01010111111: color_data = 12'b011011011110;

		11'b01011000000: color_data = 12'b011011011110;
		11'b01011000001: color_data = 12'b000000000000;
		11'b01011000010: color_data = 12'b101100100000;
		11'b01011000011: color_data = 12'b101100100000;
		11'b01011000100: color_data = 12'b101100100000;
		11'b01011000101: color_data = 12'b101100100000;
		11'b01011000110: color_data = 12'b000000000000;
		11'b01011000111: color_data = 12'b111111111111;
		11'b01011001000: color_data = 12'b101100100000;
		11'b01011001001: color_data = 12'b101100100000;
		11'b01011001010: color_data = 12'b101100100000;
		11'b01011001011: color_data = 12'b101100100000;
		11'b01011001100: color_data = 12'b000000000000;
		11'b01011001101: color_data = 12'b000000000000;
		11'b01011001110: color_data = 12'b011011011110;
		11'b01011001111: color_data = 12'b011011011110;

		11'b01011010000: color_data = 12'b011011011110;
		11'b01011010001: color_data = 12'b011011011110;
		11'b01011010010: color_data = 12'b000000000000;
		11'b01011010011: color_data = 12'b000000000000;
		11'b01011010100: color_data = 12'b101100100000;
		11'b01011010101: color_data = 12'b101100100000;
		11'b01011010110: color_data = 12'b000000000000;
		11'b01011010111: color_data = 12'b101100100000;
		11'b01011011000: color_data = 12'b101100100000;
		11'b01011011001: color_data = 12'b101100100000;
		11'b01011011010: color_data = 12'b101100100000;
		11'b01011011011: color_data = 12'b000000000000;
		11'b01011011100: color_data = 12'b000000000000;
		11'b01011011101: color_data = 12'b011011011110;
		11'b01011011110: color_data = 12'b011011011110;
		11'b01011011111: color_data = 12'b011011011110;

		11'b01011100000: color_data = 12'b011011011110;
		11'b01011100001: color_data = 12'b011011011110;
		11'b01011100010: color_data = 12'b011011011110;
		11'b01011100011: color_data = 12'b011011011110;
		11'b01011100100: color_data = 12'b000000000000;
		11'b01011100101: color_data = 12'b000000000000;
		11'b01011100110: color_data = 12'b000000000000;
		11'b01011100111: color_data = 12'b000000000000;
		11'b01011101000: color_data = 12'b000000000000;
		11'b01011101001: color_data = 12'b000000000000;
		11'b01011101010: color_data = 12'b000000000000;
		11'b01011101011: color_data = 12'b000000000000;
		11'b01011101100: color_data = 12'b011011011110;
		11'b01011101101: color_data = 12'b011011011110;
		11'b01011101110: color_data = 12'b011011011110;
		11'b01011101111: color_data = 12'b011011011110;

		11'b01011110000: color_data = 12'b011011011110;
		11'b01011110001: color_data = 12'b011011011110;
		11'b01011110010: color_data = 12'b011011011110;
		11'b01011110011: color_data = 12'b011011011110;
		11'b01011110100: color_data = 12'b011011011110;
		11'b01011110101: color_data = 12'b011011011110;
		11'b01011110110: color_data = 12'b011011011110;
		11'b01011110111: color_data = 12'b011011011110;
		11'b01011111000: color_data = 12'b011011011110;
		11'b01011111001: color_data = 12'b011011011110;
		11'b01011111010: color_data = 12'b011011011110;
		11'b01011111011: color_data = 12'b011011011110;
		11'b01011111100: color_data = 12'b011011011110;
		11'b01011111101: color_data = 12'b011011011110;
		11'b01011111110: color_data = 12'b011011011110;
		11'b01011111111: color_data = 12'b011011011110;

		11'b01100000000: color_data = 12'b000000000000;
		11'b01100000001: color_data = 12'b111111111111;
		11'b01100000010: color_data = 12'b000010110000;
		11'b01100000011: color_data = 12'b000001110000;
		11'b01100000100: color_data = 12'b000000000000;
		11'b01100000101: color_data = 12'b000000000000;
		11'b01100000110: color_data = 12'b011011011110;
		11'b01100000111: color_data = 12'b000000000000;
		11'b01100001000: color_data = 12'b000000000000;
		11'b01100001001: color_data = 12'b000000000000;
		11'b01100001010: color_data = 12'b000000000000;
		11'b01100001011: color_data = 12'b011011011110;
		11'b01100001100: color_data = 12'b000000000000;
		11'b01100001101: color_data = 12'b000000000000;
		11'b01100001110: color_data = 12'b011011011110;
		11'b01100001111: color_data = 12'b011011011110;

		11'b01100010000: color_data = 12'b000000000000;
		11'b01100010001: color_data = 12'b111111111111;
		11'b01100010010: color_data = 12'b000011110000;
		11'b01100010011: color_data = 12'b000010110000;
		11'b01100010100: color_data = 12'b000000000000;
		11'b01100010101: color_data = 12'b111111111111;
		11'b01100010110: color_data = 12'b000000000000;
		11'b01100010111: color_data = 12'b111111111111;
		11'b01100011000: color_data = 12'b111110000000;
		11'b01100011001: color_data = 12'b111110000000;
		11'b01100011010: color_data = 12'b101100100000;
		11'b01100011011: color_data = 12'b000000000000;
		11'b01100011100: color_data = 12'b111111111111;
		11'b01100011101: color_data = 12'b000000000000;
		11'b01100011110: color_data = 12'b000000000000;
		11'b01100011111: color_data = 12'b000000000000;

		11'b01100100000: color_data = 12'b000000000000;
		11'b01100100001: color_data = 12'b111111111111;
		11'b01100100010: color_data = 12'b000011110000;
		11'b01100100011: color_data = 12'b000010110000;
		11'b01100100100: color_data = 12'b000000000000;
		11'b01100100101: color_data = 12'b111111111111;
		11'b01100100110: color_data = 12'b000000000000;
		11'b01100100111: color_data = 12'b111110000000;
		11'b01100101000: color_data = 12'b101100100000;
		11'b01100101001: color_data = 12'b101100100000;
		11'b01100101010: color_data = 12'b101100100000;
		11'b01100101011: color_data = 12'b000000000000;
		11'b01100101100: color_data = 12'b111111111111;
		11'b01100101101: color_data = 12'b000000000000;
		11'b01100101110: color_data = 12'b000010110000;
		11'b01100101111: color_data = 12'b000000000000;

		11'b01100110000: color_data = 12'b000000000000;
		11'b01100110001: color_data = 12'b111111111111;
		11'b01100110010: color_data = 12'b000011110000;
		11'b01100110011: color_data = 12'b000011110000;
		11'b01100110100: color_data = 12'b000010110000;
		11'b01100110101: color_data = 12'b000000000000;
		11'b01100110110: color_data = 12'b111111111111;
		11'b01100110111: color_data = 12'b000000000000;
		11'b01100111000: color_data = 12'b000000000000;
		11'b01100111001: color_data = 12'b000000000000;
		11'b01100111010: color_data = 12'b000000000000;
		11'b01100111011: color_data = 12'b111111111111;
		11'b01100111100: color_data = 12'b000000000000;
		11'b01100111101: color_data = 12'b000010110000;
		11'b01100111110: color_data = 12'b000000000000;
		11'b01100111111: color_data = 12'b011011011110;

		11'b01101000000: color_data = 12'b011011011110;
		11'b01101000001: color_data = 12'b000000000000;
		11'b01101000010: color_data = 12'b000000000000;
		11'b01101000011: color_data = 12'b000000000000;
		11'b01101000100: color_data = 12'b000010110000;
		11'b01101000101: color_data = 12'b000000000000;
		11'b01101000110: color_data = 12'b000000000000;
		11'b01101000111: color_data = 12'b111111111111;
		11'b01101001000: color_data = 12'b111111111111;
		11'b01101001001: color_data = 12'b111111111111;
		11'b01101001010: color_data = 12'b111111111111;
		11'b01101001011: color_data = 12'b111111111111;
		11'b01101001100: color_data = 12'b000000000000;
		11'b01101001101: color_data = 12'b000010110000;
		11'b01101001110: color_data = 12'b000000000000;
		11'b01101001111: color_data = 12'b011011011110;

		11'b01101010000: color_data = 12'b000000000000;
		11'b01101010001: color_data = 12'b111110000000;
		11'b01101010010: color_data = 12'b111110000000;
		11'b01101010011: color_data = 12'b111110000000;
		11'b01101010100: color_data = 12'b000000000000;
		11'b01101010101: color_data = 12'b111110000000;
		11'b01101010110: color_data = 12'b111110000000;
		11'b01101010111: color_data = 12'b000000000000;
		11'b01101011000: color_data = 12'b000000000000;
		11'b01101011001: color_data = 12'b000000000000;
		11'b01101011010: color_data = 12'b000000000000;
		11'b01101011011: color_data = 12'b000000000000;
		11'b01101011100: color_data = 12'b000010110000;
		11'b01101011101: color_data = 12'b111111111111;
		11'b01101011110: color_data = 12'b000000000000;
		11'b01101011111: color_data = 12'b011011011110;

		11'b01101100000: color_data = 12'b000000000000;
		11'b01101100001: color_data = 12'b111110000000;
		11'b01101100010: color_data = 12'b111110000000;
		11'b01101100011: color_data = 12'b111110000000;
		11'b01101100100: color_data = 12'b111110000000;
		11'b01101100101: color_data = 12'b111110000000;
		11'b01101100110: color_data = 12'b000000000000;
		11'b01101100111: color_data = 12'b000010110000;
		11'b01101101000: color_data = 12'b000010110000;
		11'b01101101001: color_data = 12'b000010110000;
		11'b01101101010: color_data = 12'b000010110000;
		11'b01101101011: color_data = 12'b000010110000;
		11'b01101101100: color_data = 12'b111111111111;
		11'b01101101101: color_data = 12'b000000000000;
		11'b01101101110: color_data = 12'b011011011110;
		11'b01101101111: color_data = 12'b011011011110;

		11'b01101110000: color_data = 12'b000000000000;
		11'b01101110001: color_data = 12'b111110000000;
		11'b01101110010: color_data = 12'b111110000000;
		11'b01101110011: color_data = 12'b111110000000;
		11'b01101110100: color_data = 12'b000000000000;
		11'b01101110101: color_data = 12'b000000000000;
		11'b01101110110: color_data = 12'b111111111111;
		11'b01101110111: color_data = 12'b111111111111;
		11'b01101111000: color_data = 12'b111111111111;
		11'b01101111001: color_data = 12'b000000000000;
		11'b01101111010: color_data = 12'b000000000000;
		11'b01101111011: color_data = 12'b111111111111;
		11'b01101111100: color_data = 12'b111111111111;
		11'b01101111101: color_data = 12'b000000000000;
		11'b01101111110: color_data = 12'b011011011110;
		11'b01101111111: color_data = 12'b011011011110;

		11'b01110000000: color_data = 12'b011011011110;
		11'b01110000001: color_data = 12'b000000000000;
		11'b01110000010: color_data = 12'b000000000000;
		11'b01110000011: color_data = 12'b000000000000;
		11'b01110000100: color_data = 12'b111111111111;
		11'b01110000101: color_data = 12'b111111111111;
		11'b01110000110: color_data = 12'b111111111111;
		11'b01110000111: color_data = 12'b111111111111;
		11'b01110001000: color_data = 12'b000000000000;
		11'b01110001001: color_data = 12'b000010110000;
		11'b01110001010: color_data = 12'b000011110000;
		11'b01110001011: color_data = 12'b000000000000;
		11'b01110001100: color_data = 12'b000000000000;
		11'b01110001101: color_data = 12'b000000000000;
		11'b01110001110: color_data = 12'b011011011110;
		11'b01110001111: color_data = 12'b011011011110;

		11'b01110010000: color_data = 12'b000000000000;
		11'b01110010001: color_data = 12'b000000000000;
		11'b01110010010: color_data = 12'b000000000000;
		11'b01110010011: color_data = 12'b111111111111;
		11'b01110010100: color_data = 12'b111111111111;
		11'b01110010101: color_data = 12'b111111111111;
		11'b01110010110: color_data = 12'b111111111111;
		11'b01110010111: color_data = 12'b111111111111;
		11'b01110011000: color_data = 12'b000000000000;
		11'b01110011001: color_data = 12'b000010110000;
		11'b01110011010: color_data = 12'b000000000000;
		11'b01110011011: color_data = 12'b101100100000;
		11'b01110011100: color_data = 12'b101100100000;
		11'b01110011101: color_data = 12'b101100100000;
		11'b01110011110: color_data = 12'b000000000000;
		11'b01110011111: color_data = 12'b011011011110;

		11'b01110100000: color_data = 12'b000000000000;
		11'b01110100001: color_data = 12'b111111111111;
		11'b01110100010: color_data = 12'b101100100000;
		11'b01110100011: color_data = 12'b000000000000;
		11'b01110100100: color_data = 12'b000000000000;
		11'b01110100101: color_data = 12'b111111111111;
		11'b01110100110: color_data = 12'b111111111111;
		11'b01110100111: color_data = 12'b111111111111;
		11'b01110101000: color_data = 12'b000000000000;
		11'b01110101001: color_data = 12'b000000000000;
		11'b01110101010: color_data = 12'b101100100000;
		11'b01110101011: color_data = 12'b101100100000;
		11'b01110101100: color_data = 12'b101100100000;
		11'b01110101101: color_data = 12'b101100100000;
		11'b01110101110: color_data = 12'b101100100000;
		11'b01110101111: color_data = 12'b000000000000;

		11'b01110110000: color_data = 12'b000000000000;
		11'b01110110001: color_data = 12'b101100100000;
		11'b01110110010: color_data = 12'b101100100000;
		11'b01110110011: color_data = 12'b101100100000;
		11'b01110110100: color_data = 12'b101100100000;
		11'b01110110101: color_data = 12'b000000000000;
		11'b01110110110: color_data = 12'b000000000000;
		11'b01110110111: color_data = 12'b000000000000;
		11'b01110111000: color_data = 12'b000000000000;
		11'b01110111001: color_data = 12'b000000000000;
		11'b01110111010: color_data = 12'b101100100000;
		11'b01110111011: color_data = 12'b101100100000;
		11'b01110111100: color_data = 12'b101100100000;
		11'b01110111101: color_data = 12'b101100100000;
		11'b01110111110: color_data = 12'b000000000000;
		11'b01110111111: color_data = 12'b011011011110;

		11'b01111000000: color_data = 12'b011011011110;
		11'b01111000001: color_data = 12'b000000000000;
		11'b01111000010: color_data = 12'b101100100000;
		11'b01111000011: color_data = 12'b101100100000;
		11'b01111000100: color_data = 12'b101100100000;
		11'b01111000101: color_data = 12'b101100100000;
		11'b01111000110: color_data = 12'b101100100000;
		11'b01111000111: color_data = 12'b000000000000;
		11'b01111001000: color_data = 12'b000000000000;
		11'b01111001001: color_data = 12'b111111111111;
		11'b01111001010: color_data = 12'b101100100000;
		11'b01111001011: color_data = 12'b101100100000;
		11'b01111001100: color_data = 12'b101100100000;
		11'b01111001101: color_data = 12'b000000000000;
		11'b01111001110: color_data = 12'b011011011110;
		11'b01111001111: color_data = 12'b011011011110;

		11'b01111010000: color_data = 12'b011011011110;
		11'b01111010001: color_data = 12'b011011011110;
		11'b01111010010: color_data = 12'b000000000000;
		11'b01111010011: color_data = 12'b101100100000;
		11'b01111010100: color_data = 12'b101100100000;
		11'b01111010101: color_data = 12'b101100100000;
		11'b01111010110: color_data = 12'b000000000000;
		11'b01111010111: color_data = 12'b011011011110;
		11'b01111011000: color_data = 12'b000000000000;
		11'b01111011001: color_data = 12'b101100100000;
		11'b01111011010: color_data = 12'b101100100000;
		11'b01111011011: color_data = 12'b101100100000;
		11'b01111011100: color_data = 12'b000000000000;
		11'b01111011101: color_data = 12'b011011011110;
		11'b01111011110: color_data = 12'b011011011110;
		11'b01111011111: color_data = 12'b011011011110;

		11'b01111100000: color_data = 12'b011011011110;
		11'b01111100001: color_data = 12'b011011011110;
		11'b01111100010: color_data = 12'b011011011110;
		11'b01111100011: color_data = 12'b000000000000;
		11'b01111100100: color_data = 12'b000000000000;
		11'b01111100101: color_data = 12'b000000000000;
		11'b01111100110: color_data = 12'b011011011110;
		11'b01111100111: color_data = 12'b011011011110;
		11'b01111101000: color_data = 12'b000000000000;
		11'b01111101001: color_data = 12'b000000000000;
		11'b01111101010: color_data = 12'b000000000000;
		11'b01111101011: color_data = 12'b000000000000;
		11'b01111101100: color_data = 12'b011011011110;
		11'b01111101101: color_data = 12'b011011011110;
		11'b01111101110: color_data = 12'b011011011110;
		11'b01111101111: color_data = 12'b011011011110;

		11'b01111110000: color_data = 12'b011011011110;
		11'b01111110001: color_data = 12'b011011011110;
		11'b01111110010: color_data = 12'b011011011110;
		11'b01111110011: color_data = 12'b011011011110;
		11'b01111110100: color_data = 12'b011011011110;
		11'b01111110101: color_data = 12'b011011011110;
		11'b01111110110: color_data = 12'b011011011110;
		11'b01111110111: color_data = 12'b011011011110;
		11'b01111111000: color_data = 12'b011011011110;
		11'b01111111001: color_data = 12'b011011011110;
		11'b01111111010: color_data = 12'b011011011110;
		11'b01111111011: color_data = 12'b011011011110;
		11'b01111111100: color_data = 12'b011011011110;
		11'b01111111101: color_data = 12'b011011011110;
		11'b01111111110: color_data = 12'b011011011110;
		11'b01111111111: color_data = 12'b011011011110;

		11'b10000000000: color_data = 12'b000000000000;
		11'b10000000001: color_data = 12'b111111111111;
		11'b10000000010: color_data = 12'b000011110000;
		11'b10000000011: color_data = 12'b000001110000;
		11'b10000000100: color_data = 12'b000000000000;
		11'b10000000101: color_data = 12'b000000000000;
		11'b10000000110: color_data = 12'b011011011110;
		11'b10000000111: color_data = 12'b000000000000;
		11'b10000001000: color_data = 12'b000000000000;
		11'b10000001001: color_data = 12'b000000000000;
		11'b10000001010: color_data = 12'b000000000000;
		11'b10000001011: color_data = 12'b011011011110;
		11'b10000001100: color_data = 12'b000000000000;
		11'b10000001101: color_data = 12'b000000000000;
		11'b10000001110: color_data = 12'b011011011110;
		11'b10000001111: color_data = 12'b011011011110;

		11'b10000010000: color_data = 12'b000000000000;
		11'b10000010001: color_data = 12'b111111111111;
		11'b10000010010: color_data = 12'b111111111111;
		11'b10000010011: color_data = 12'b000011110000;
		11'b10000010100: color_data = 12'b000000000000;
		11'b10000010101: color_data = 12'b111111111111;
		11'b10000010110: color_data = 12'b000000000000;
		11'b10000010111: color_data = 12'b111111111111;
		11'b10000011000: color_data = 12'b111110000000;
		11'b10000011001: color_data = 12'b111110000000;
		11'b10000011010: color_data = 12'b101100100000;
		11'b10000011011: color_data = 12'b000000000000;
		11'b10000011100: color_data = 12'b111111111111;
		11'b10000011101: color_data = 12'b000000000000;
		11'b10000011110: color_data = 12'b000000000000;
		11'b10000011111: color_data = 12'b000000000000;

		11'b10000100000: color_data = 12'b000000000000;
		11'b10000100001: color_data = 12'b111111111111;
		11'b10000100010: color_data = 12'b111111111111;
		11'b10000100011: color_data = 12'b111111111111;
		11'b10000100100: color_data = 12'b000000000000;
		11'b10000100101: color_data = 12'b111111111111;
		11'b10000100110: color_data = 12'b000000000000;
		11'b10000100111: color_data = 12'b111110000000;
		11'b10000101000: color_data = 12'b101100100000;
		11'b10000101001: color_data = 12'b101100100000;
		11'b10000101010: color_data = 12'b101100100000;
		11'b10000101011: color_data = 12'b000000000000;
		11'b10000101100: color_data = 12'b111111111111;
		11'b10000101101: color_data = 12'b000000000000;
		11'b10000101110: color_data = 12'b000010110000;
		11'b10000101111: color_data = 12'b000000000000;

		11'b10000110000: color_data = 12'b000000000000;
		11'b10000110001: color_data = 12'b111111111111;
		11'b10000110010: color_data = 12'b111111111111;
		11'b10000110011: color_data = 12'b111111111111;
		11'b10000110100: color_data = 12'b111111111111;
		11'b10000110101: color_data = 12'b000000000000;
		11'b10000110110: color_data = 12'b111111111111;
		11'b10000110111: color_data = 12'b000000000000;
		11'b10000111000: color_data = 12'b000000000000;
		11'b10000111001: color_data = 12'b000000000000;
		11'b10000111010: color_data = 12'b000000000000;
		11'b10000111011: color_data = 12'b111111111111;
		11'b10000111100: color_data = 12'b000000000000;
		11'b10000111101: color_data = 12'b111111111111;
		11'b10000111110: color_data = 12'b000000000000;
		11'b10000111111: color_data = 12'b011011011110;

		11'b10001000000: color_data = 12'b000000000000;
		11'b10001000001: color_data = 12'b111111111111;
		11'b10001000010: color_data = 12'b111111111111;
		11'b10001000011: color_data = 12'b111111111111;
		11'b10001000100: color_data = 12'b000000000000;
		11'b10001000101: color_data = 12'b000000000000;
		11'b10001000110: color_data = 12'b000000000000;
		11'b10001000111: color_data = 12'b111111111111;
		11'b10001001000: color_data = 12'b111111111111;
		11'b10001001001: color_data = 12'b111111111111;
		11'b10001001010: color_data = 12'b111111111111;
		11'b10001001011: color_data = 12'b111111111111;
		11'b10001001100: color_data = 12'b000000000000;
		11'b10001001101: color_data = 12'b111111111111;
		11'b10001001110: color_data = 12'b000000000000;
		11'b10001001111: color_data = 12'b011011011110;

		11'b10001010000: color_data = 12'b011011011110;
		11'b10001010001: color_data = 12'b000000000000;
		11'b10001010010: color_data = 12'b111111111111;
		11'b10001010011: color_data = 12'b111111111111;
		11'b10001010100: color_data = 12'b000000000000;
		11'b10001010101: color_data = 12'b111110000000;
		11'b10001010110: color_data = 12'b111110000000;
		11'b10001010111: color_data = 12'b000000000000;
		11'b10001011000: color_data = 12'b000000000000;
		11'b10001011001: color_data = 12'b000000000000;
		11'b10001011010: color_data = 12'b000000000000;
		11'b10001011011: color_data = 12'b000000000000;
		11'b10001011100: color_data = 12'b111111111111;
		11'b10001011101: color_data = 12'b111111111111;
		11'b10001011110: color_data = 12'b000000000000;
		11'b10001011111: color_data = 12'b011011011110;

		11'b10001100000: color_data = 12'b011011011110;
		11'b10001100001: color_data = 12'b000000000000;
		11'b10001100010: color_data = 12'b111111111111;
		11'b10001100011: color_data = 12'b111111111111;
		11'b10001100100: color_data = 12'b111111111111;
		11'b10001100101: color_data = 12'b000000000000;
		11'b10001100110: color_data = 12'b111110000000;
		11'b10001100111: color_data = 12'b111110000000;
		11'b10001101000: color_data = 12'b000000000000;
		11'b10001101001: color_data = 12'b111111111111;
		11'b10001101010: color_data = 12'b111111111111;
		11'b10001101011: color_data = 12'b111111111111;
		11'b10001101100: color_data = 12'b111111111111;
		11'b10001101101: color_data = 12'b000000000000;
		11'b10001101110: color_data = 12'b011011011110;
		11'b10001101111: color_data = 12'b011011011110;

		11'b10001110000: color_data = 12'b011011011110;
		11'b10001110001: color_data = 12'b011011011110;
		11'b10001110010: color_data = 12'b000000000000;
		11'b10001110011: color_data = 12'b111111111111;
		11'b10001110100: color_data = 12'b111111111111;
		11'b10001110101: color_data = 12'b111111111111;
		11'b10001110110: color_data = 12'b000000000000;
		11'b10001110111: color_data = 12'b111110000000;
		11'b10001111000: color_data = 12'b000000000000;
		11'b10001111001: color_data = 12'b111111111111;
		11'b10001111010: color_data = 12'b111111111111;
		11'b10001111011: color_data = 12'b111111111111;
		11'b10001111100: color_data = 12'b111111111111;
		11'b10001111101: color_data = 12'b000000000000;
		11'b10001111110: color_data = 12'b011011011110;
		11'b10001111111: color_data = 12'b011011011110;

		11'b10010000000: color_data = 12'b011011011110;
		11'b10010000001: color_data = 12'b011011011110;
		11'b10010000010: color_data = 12'b000000000000;
		11'b10010000011: color_data = 12'b111111111111;
		11'b10010000100: color_data = 12'b111111111111;
		11'b10010000101: color_data = 12'b000000000000;
		11'b10010000110: color_data = 12'b111110000000;
		11'b10010000111: color_data = 12'b111110000000;
		11'b10010001000: color_data = 12'b111110000000;
		11'b10010001001: color_data = 12'b000000000000;
		11'b10010001010: color_data = 12'b000000000000;
		11'b10010001011: color_data = 12'b000000000000;
		11'b10010001100: color_data = 12'b000000000000;
		11'b10010001101: color_data = 12'b000000000000;
		11'b10010001110: color_data = 12'b011011011110;
		11'b10010001111: color_data = 12'b011011011110;

		11'b10010010000: color_data = 12'b011011011110;
		11'b10010010001: color_data = 12'b011011011110;
		11'b10010010010: color_data = 12'b011011011110;
		11'b10010010011: color_data = 12'b000000000000;
		11'b10010010100: color_data = 12'b111111111111;
		11'b10010010101: color_data = 12'b000000000000;
		11'b10010010110: color_data = 12'b111110000000;
		11'b10010010111: color_data = 12'b111110000000;
		11'b10010011000: color_data = 12'b111110000000;
		11'b10010011001: color_data = 12'b000000000000;
		11'b10010011010: color_data = 12'b101100100000;
		11'b10010011011: color_data = 12'b101100100000;
		11'b10010011100: color_data = 12'b101100100000;
		11'b10010011101: color_data = 12'b000000000000;
		11'b10010011110: color_data = 12'b011011011110;
		11'b10010011111: color_data = 12'b011011011110;

		11'b10010100000: color_data = 12'b011011011110;
		11'b10010100001: color_data = 12'b011011011110;
		11'b10010100010: color_data = 12'b011011011110;
		11'b10010100011: color_data = 12'b011011011110;
		11'b10010100100: color_data = 12'b000000000000;
		11'b10010100101: color_data = 12'b111111111111;
		11'b10010100110: color_data = 12'b000000000000;
		11'b10010100111: color_data = 12'b000000000000;
		11'b10010101000: color_data = 12'b000000000000;
		11'b10010101001: color_data = 12'b000000000000;
		11'b10010101010: color_data = 12'b101100100000;
		11'b10010101011: color_data = 12'b101100100000;
		11'b10010101100: color_data = 12'b101100100000;
		11'b10010101101: color_data = 12'b000000000000;
		11'b10010101110: color_data = 12'b011011011110;
		11'b10010101111: color_data = 12'b011011011110;

		11'b10010110000: color_data = 12'b011011011110;
		11'b10010110001: color_data = 12'b011011011110;
		11'b10010110010: color_data = 12'b011011011110;
		11'b10010110011: color_data = 12'b011011011110;
		11'b10010110100: color_data = 12'b011011011110;
		11'b10010110101: color_data = 12'b000000000000;
		11'b10010110110: color_data = 12'b000000000000;
		11'b10010110111: color_data = 12'b000010110000;
		11'b10010111000: color_data = 12'b111111111111;
		11'b10010111001: color_data = 12'b000000000000;
		11'b10010111010: color_data = 12'b101100100000;
		11'b10010111011: color_data = 12'b101100100000;
		11'b10010111100: color_data = 12'b101100100000;
		11'b10010111101: color_data = 12'b000000000000;
		11'b10010111110: color_data = 12'b011011011110;
		11'b10010111111: color_data = 12'b011011011110;

		11'b10011000000: color_data = 12'b011011011110;
		11'b10011000001: color_data = 12'b011011011110;
		11'b10011000010: color_data = 12'b011011011110;
		11'b10011000011: color_data = 12'b011011011110;
		11'b10011000100: color_data = 12'b011011011110;
		11'b10011000101: color_data = 12'b011011011110;
		11'b10011000110: color_data = 12'b011011011110;
		11'b10011000111: color_data = 12'b000000000000;
		11'b10011001000: color_data = 12'b000010110000;
		11'b10011001001: color_data = 12'b000000000000;
		11'b10011001010: color_data = 12'b101100100000;
		11'b10011001011: color_data = 12'b101100100000;
		11'b10011001100: color_data = 12'b101100100000;
		11'b10011001101: color_data = 12'b000000000000;
		11'b10011001110: color_data = 12'b011011011110;
		11'b10011001111: color_data = 12'b011011011110;

		11'b10011010000: color_data = 12'b011011011110;
		11'b10011010001: color_data = 12'b011011011110;
		11'b10011010010: color_data = 12'b011011011110;
		11'b10011010011: color_data = 12'b011011011110;
		11'b10011010100: color_data = 12'b011011011110;
		11'b10011010101: color_data = 12'b011011011110;
		11'b10011010110: color_data = 12'b011011011110;
		11'b10011010111: color_data = 12'b011011011110;
		11'b10011011000: color_data = 12'b000000000000;
		11'b10011011001: color_data = 12'b000000000000;
		11'b10011011010: color_data = 12'b101100100000;
		11'b10011011011: color_data = 12'b101100100000;
		11'b10011011100: color_data = 12'b101100100000;
		11'b10011011101: color_data = 12'b000000000000;
		11'b10011011110: color_data = 12'b011011011110;
		11'b10011011111: color_data = 12'b011011011110;

		11'b10011100000: color_data = 12'b011011011110;
		11'b10011100001: color_data = 12'b011011011110;
		11'b10011100010: color_data = 12'b011011011110;
		11'b10011100011: color_data = 12'b011011011110;
		11'b10011100100: color_data = 12'b011011011110;
		11'b10011100101: color_data = 12'b011011011110;
		11'b10011100110: color_data = 12'b011011011110;
		11'b10011100111: color_data = 12'b011011011110;
		11'b10011101000: color_data = 12'b011011011110;
		11'b10011101001: color_data = 12'b011011011110;
		11'b10011101010: color_data = 12'b000000000000;
		11'b10011101011: color_data = 12'b111111111111;
		11'b10011101100: color_data = 12'b101100100000;
		11'b10011101101: color_data = 12'b000000000000;
		11'b10011101110: color_data = 12'b011011011110;
		11'b10011101111: color_data = 12'b011011011110;

		11'b10011110000: color_data = 12'b011011011110;
		11'b10011110001: color_data = 12'b011011011110;
		11'b10011110010: color_data = 12'b011011011110;
		11'b10011110011: color_data = 12'b011011011110;
		11'b10011110100: color_data = 12'b011011011110;
		11'b10011110101: color_data = 12'b011011011110;
		11'b10011110110: color_data = 12'b011011011110;
		11'b10011110111: color_data = 12'b011011011110;
		11'b10011111000: color_data = 12'b011011011110;
		11'b10011111001: color_data = 12'b011011011110;
		11'b10011111010: color_data = 12'b011011011110;
		11'b10011111011: color_data = 12'b000000000000;
		11'b10011111100: color_data = 12'b000000000000;
		11'b10011111101: color_data = 12'b000000000000;
		11'b10011111110: color_data = 12'b011011011110;
		11'b10011111111: color_data = 12'b011011011110;

		default: color_data = 12'b000000000000;
	endcase
endmodule